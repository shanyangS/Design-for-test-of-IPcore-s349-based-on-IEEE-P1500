module sel_gen
(
	input wby_shift,wir_wpc,wir_extest,wir_intest,
	output[3:0] sel_o,
);

always@(*)
	if(wby_shift = 1)

endmodule
